`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   08:38:00 09/04/2023
// Design Name:   cpu_checker
// Module Name:   /home/co-eda/ISE/T-1109-397/tb_cpu_checker.v
// Project Name:  T-1109-397
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: cpu_checker
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module tb_cpu_checker;

	// Inputs
	reg clk;
	reg reset;
	reg [7:0] char;
	reg [15:0] freq;
	reg finish;

	// Outputs
	wire [1:0] format_type;
	wire [3:0] error_code;

	// debug
	// wire [3:0] status_output;
	// wire [3:0] error_output;
	// wire [31:0] pc_store_output;
	// wire [31:0] addr_store_output;

	// Instantiate the Unit Under Test (UUT)
	cpu_checker uut (
		.clk(clk), 
		.reset(reset), 
		.char(char), 
		.freq(freq), 
		.format_type(format_type), 
		.error_code(error_code)
		// debug
		// .status_output(status_output),
		// .error_output(error_output),
		// .pc_store_output(pc_store_output),
		// .addr_store_output(addr_store_output)
	);

	always @(posedge clk) begin
		if (!reset && !finish) begin
			$display("%d %d", format_type, error_code);
		end
	end

	initial begin
		// Initialize Inputs
		clk = 0;
		reset = 1;
		char = 0;
		freq = 4;
		finish = 0;

		#10 reset = 0;
		#2 char = "^";
		#2 char = "2";
		#2 char = "4";
		#2 char = "2";
		#2 char = "@";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "3";
		#2 char = "0";
		#2 char = "f";
		#2 char = "4";
		#2 char = ":";
		#2 char = " ";
		#2 char = "$";
		#2 char = "3";
		#2 char = "1";
		#2 char = " ";
		#2 char = "<";
		#2 char = "=";
		#2 char = "1";
		#2 char = "2";
		#2 char = "3";
		#2 char = "4";
		#2 char = "5";
		#2 char = "6";
		#2 char = "7";
		#2 char = "8";
		#2 char = "#";
		#2 char = "^";
		#2 char = "2";
		#2 char = "4";
		#2 char = "2";
		#2 char = "@";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "3";
		#2 char = "0";
		#2 char = "f";
		#2 char = "4";
		#2 char = ":";
		#2 char = " ";
		#2 char = "$";
		#2 char = "3";
		#2 char = "1";
		#2 char = " ";
		#2 char = "<";
		#2 char = "=";
		#2 char = "1";
		#2 char = "2";
		#2 char = "3";
		#2 char = "2";
		#2 char = "1";
		#2 char = "5";
		#2 char = "#";
		#2 char = "^";
		#2 char = "2";
		#2 char = "4";
		#2 char = "2";
		#2 char = "@";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "3";
		#2 char = "0";
		#2 char = "f";
		#2 char = "4";
		#2 char = ":";
		#2 char = " ";
		#2 char = "$";
		#2 char = "3";
		#2 char = "1";
		#2 char = " ";
		#2 char = "<";
		#2 char = "=";
		#2 char = "1";
		#2 char = "2";
		#2 char = "3";
		#2 char = "2";
		#2 char = "1";
		#2 char = "5";
		#2 char = "8";
		#2 char = "9";
		#2 char = "9";
		#2 char = "8";
		#2 char = "#";
		#2 char = "^";
		#2 char = "2";
		#2 char = "4";
		#2 char = "2";
		#2 char = "@";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "3";
		#2 char = "0";
		#2 char = "f";
		#2 char = "4";
		#2 char = ":";
		#2 char = " ";
		#2 char = "$";
		#2 char = "3";
		#2 char = "1";
		#2 char = " ";
		#2 char = "<";
		#2 char = "=";
		#2 char = "#";
		#2 char = "^";
		#2 char = "2";
		#2 char = "4";
		#2 char = "2";
		#2 char = "@";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "3";
		#2 char = "0";
		#2 char = "f";
		#2 char = "4";
		#2 char = ":";
		#2 char = " ";
		#2 char = "$";
		#2 char = "3";
		#2 char = "1";
		#2 char = " ";
		#2 char = "<";
		#2 char = "=";
		#2 char = " ";
		#2 char = " ";
		#2 char = " ";
		#2 char = "1";
		#2 char = "2";
		#2 char = "3";
		#2 char = "2";
		#2 char = "1";
		#2 char = "5";
		#2 char = " ";
		#2 char = "#";
		#2 char = "^";
		#2 char = "2";
		#2 char = "4";
		#2 char = "2";
		#2 char = "@";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "3";
		#2 char = "0";
		#2 char = "f";
		#2 char = "4";
		#2 char = ":";
		#2 char = " ";
		#2 char = "$";
		#2 char = "3";
		#2 char = "1";
		#2 char = " ";
		#2 char = "<";
		#2 char = "=";
		#2 char = " ";
		#2 char = " ";
		#2 char = " ";
		#2 char = "a";
		#2 char = "b";
		#2 char = "1";
		#2 char = "2";
		#2 char = "3";
		#2 char = "2";
		#2 char = "1";
		#2 char = "5";
		#2 char = " ";
		#2 char = "#";
		#2 char = "^";
		#2 char = "2";
		#2 char = "4";
		#2 char = "2";
		#2 char = "@";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "3";
		#2 char = "0";
		#2 char = "f";
		#2 char = "4";
		#2 char = ":";
		#2 char = " ";
		#2 char = "$";
		#2 char = "3";
		#2 char = "1";
		#2 char = " ";
		#2 char = "<";
		#2 char = "=";
		#2 char = " ";
		#2 char = " ";
		#2 char = " ";
		#2 char = "A";
		#2 char = "b";
		#2 char = "1";
		#2 char = "2";
		#2 char = "3";
		#2 char = "2";
		#2 char = "1";
		#2 char = "5";
		#2 char = " ";
		#2 char = "#";
		#2 char = "^";
		#2 char = "3";
		#2 char = "3";
		#2 char = "8";
		#2 char = "@";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "3";
		#2 char = "1";
		#2 char = "3";
		#2 char = "0";
		#2 char = ":";
		#2 char = " ";
		#2 char = "*";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "8";
		#2 char = "8";
		#2 char = " ";
		#2 char = "<";
		#2 char = "=";
		#2 char = " ";
		#2 char = "F";
		#2 char = "f";
		#2 char = "f";
		#2 char = "f";
		#2 char = "b";
		#2 char = "5";
		#2 char = "2";
		#2 char = "8";
		#2 char = "#";
		#2 char = "^";
		#2 char = "3";
		#2 char = "3";
		#2 char = "8";
		#2 char = "@";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "3";
		#2 char = "1";
		#2 char = "3";
		#2 char = "0";
		#2 char = ":";
		#2 char = " ";
		#2 char = "*";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "8";
		#2 char = "8";
		#2 char = " ";
		#2 char = "<";
		#2 char = "=";
		#2 char = " ";
		#2 char = "f";
		#2 char = "f";
		#2 char = "f";
		#2 char = "f";
		#2 char = "b";
		#2 char = "5";
		#2 char = "2";
		#2 char = "8";
		#2 char = "#";
		#2 char = "^";
		#2 char = "3";
		#2 char = "3";
		#2 char = "8";
		#2 char = "@";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "3";
		#2 char = "1";
		#2 char = "3";
		#2 char = "0";
		#2 char = ":";
		#2 char = " ";
		#2 char = "*";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "8";
		#2 char = "8";
		#2 char = " ";
		#2 char = "<";
		#2 char = "=";
		#2 char = "#";
		#2 char = "^";
		#2 char = "3";
		#2 char = "3";
		#2 char = "8";
		#2 char = "@";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "3";
		#2 char = "1";
		#2 char = "3";
		#2 char = "0";
		#2 char = ":";
		#2 char = " ";
		#2 char = "*";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "8";
		#2 char = "8";
		#2 char = " ";
		#2 char = "<";
		#2 char = "=";
		#2 char = " ";
		#2 char = "f";
		#2 char = "f";
		#2 char = "f";
		#2 char = "f";
		#2 char = "b";
		#2 char = "5";
		#2 char = "2";
		#2 char = "8";
		#2 char = "1";
		#2 char = "2";
		#2 char = "#";
		#2 char = "^";
		#2 char = "3";
		#2 char = "3";
		#2 char = "8";
		#2 char = "@";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "3";
		#2 char = "1";
		#2 char = "3";
		#2 char = "0";
		#2 char = ":";
		#2 char = " ";
		#2 char = "*";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "8";
		#2 char = "8";
		#2 char = " ";
		#2 char = "<";
		#2 char = "=";
		#2 char = " ";
		#2 char = "f";
		#2 char = "f";
		#2 char = "f";
		#2 char = "f";
		#2 char = "b";
		#2 char = "5";
		#2 char = "2";
		#2 char = "#";
		#2 char = "^";
		#2 char = "3";
		#2 char = "3";
		#2 char = "8";
		#2 char = "@";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "3";
		#2 char = "1";
		#2 char = "3";
		#2 char = "0";
		#2 char = ":";
		#2 char = " ";
		#2 char = "*";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "8";
		#2 char = "8";
		#2 char = " ";
		#2 char = "<";
		#2 char = "=";
		#2 char = " ";
		#2 char = "f";
		#2 char = "f";
		#2 char = "f";
		#2 char = "f";
		#2 char = "B";
		#2 char = "5";
		#2 char = "2";
		#2 char = "8";
		#2 char = "#";
		#2 char = "^";
		#2 char = "3";
		#2 char = "3";
		#2 char = "8";
		#2 char = "@";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "3";
		#2 char = "1";
		#2 char = "3";
		#2 char = "0";
		#2 char = ":";
		#2 char = " ";
		#2 char = "*";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "8";
		#2 char = "8";
		#2 char = " ";
		#2 char = "<";
		#2 char = "=";
		#2 char = " ";
		#2 char = "f";
		#2 char = "f";
		#2 char = "f";
		#2 char = "f";
		#2 char = "b";
		#2 char = "5";
		#2 char = "2";
		#2 char = "B";
		#2 char = "#";
		#2 char = "^";
		#2 char = "3";
		#2 char = "3";
		#2 char = "8";
		#2 char = "@";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "3";
		#2 char = "1";
		#2 char = "3";
		#2 char = "0";
		#2 char = ":";
		#2 char = " ";
		#2 char = "*";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "8";
		#2 char = "8";
		#2 char = " ";
		#2 char = "<";
		#2 char = "=";
		#2 char = " ";
		#2 char = "f";
		#2 char = "f";
		#2 char = "f";
		#2 char = "f";
		#2 char = "b";
		#2 char = "5";
		#2 char = "2";
		#2 char = "B";
		#2 char = "#";
		#2 char = "^";
		#2 char = "3";
		#2 char = "3";
		#2 char = "8";
		#2 char = "@";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "3";
		#2 char = "1";
		#2 char = "3";
		#2 char = "0";
		#2 char = ":";
		#2 char = " ";
		#2 char = "*";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "0";
		#2 char = "8";
		#2 char = "8";
		#2 char = " ";
		#2 char = "<";
		#2 char = "=";
		#2 char = " ";
		#2 char = "f";
		#2 char = "f";
		#2 char = "f";
		#2 char = "f";
		#2 char = "b";
		#2 char = "5";
		#2 char = "2";
		#2 char = "B";
		#2 char = " ";
		#2 char = "#";
		#20
		finish = 1;
	end

    always #1 clk = ~clk;
      
endmodule

